`ifndef SPI_DEFINES_VH
`define SPI_DEFINES_VH

`define DATA_LEN   8
`define DIV_WIDTH  8
`define CPOL       0
`define CPHA       0

`endif